library ieee;
package fixed_pkg is new ieee.fixed_generic_pkg;
